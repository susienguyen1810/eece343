//module FSM_top (input logic clk, Reset, left, right, hazard, brake,
//				    output logic LA,LB,LC,RA,RB,RC,
//					 input logic clr, output logic clk3
//					 );
//
//	FSM dut(
//	.left(left),
//	.right(right),
//	.hazard(hazard),
//	.brake(brake),
//	.LA(LA),
//	.LB(LB),
//	.LC(LC),
//	.RA(RA),
//	.RB(RB),
//	.RC(RC),
//	.clk(clk3),
//	.Reset(Reset)
//	);
//	
//	clkdiv uut(
//	.clk(clk),
//	.clr(clr),
//	.clk3(clk3)
//	);
//	
//endmodule
